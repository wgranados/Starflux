module rate_divider(enable, countdown_start, clock, reset, q);
	input enable; // enable signal given from user
	input reset; // reset signal given by user
	input clock; // clock signal given from CLOCK_50
	input [27:0]countdown_start; // value that this counter should start counting down from
	output reg [27:0]q; // output register we're outputting current count for this rate divider

	// start counting down from count_down_start all the way to 0
	always @(posedge clock)
	begin
		if(reset == 1'b1) // when clear_b is 0
			q <= countdown_start;
		else if(enable == 1'b1) // decrement q only when enable is high
			q <= (q == 0) ? countdown_start : q - 1'b1; // if we get to 0, then we loop back
	end

endmodule

